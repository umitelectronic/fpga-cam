----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:38:37 03/08/2012 
-- Design Name: 
-- Module Name:    block3X3 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library WORK ;
use WORK.CAMERA.ALL ;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity block3X3v2 is
		generic(LINE_SIZE : natural := 640);
		port(
			clk : in std_logic; 
			arazb : in std_logic; 
			pixel_clock, hsync, vsync : in std_logic; 
			pixel_data_in : in std_logic_vector(7 downto 0 ); 
			new_block : out std_logic ;
			block_out : out mat3);
end block3X3v2;

architecture Behavioral of block3X3v2 is
type read_pixel_state is (LOAD_VALUES1, LOAD_VALUES2, WAIT_PIXEL, END_PIXEL, END_HSYNC);
type hsync_state is	(WAIT_HSYNC, END_HSYNC);


signal pixel_state : read_pixel_state ;
signal hsync_state0 : hsync_state ;

signal block3x3 : mat3 := (((others => '0'), (others => '0'), (others => '0')), 
									((others => '0'), (others => '0'), (others => '0')), 
									((others => '0'), (others => '0'), (others => '0')));

signal k02, k12 :	signed(8 downto 0) := (others => '0');


signal line_wr, nclk: std_logic ;


signal LINE1_INPUT, LINE1_OUTPUT, LINE2_INPUT, LINE2_OUTPUT : std_logic_vector(7 downto 0) := X"00";
signal final_res : signed(31 downto 0);
signal nb_line : std_logic_vector(3 downto 0) := (others => '0');
signal pixel_counter : std_logic_vector(9 downto 0) ;
begin

nclk <= NOT clk ;

line1: ram_Nx8
	generic map(N => LINE_SIZE + 2, A => 10)
	port map(
 		clk => nclk, 
 		we => line_wr, en => '1' ,
 		do => LINE1_OUTPUT,
 		di => LINE1_INPUT,
 		addr => pixel_counter
	); 

line2: ram_Nx8
	generic map(N => LINE_SIZE + 2, A => 10)
	port map(
 		clk => nclk, 
 		we => line_wr, en => '1' ,
 		do => LINE2_OUTPUT,
 		di => LINE2_INPUT,
 		addr => pixel_counter
	); 


-- actualize matrix with values
process(clk, arazb)
begin
if arazb = '0' then 
	block3x3(0)(0) <= (others => '0') ;
	block3x3(0)(1) <= (others => '0') ; -- zeroing matrix
	block3x3(0)(2) <= (others => '0') ;
	
	block3x3(1)(0) <= (others => '0') ;
	block3x3(1)(1) <= (others => '0') ;
	block3x3(1)(2) <= (others => '0') ;
	
	block3x3(2)(0) <= (others => '0') ;
	block3x3(2)(1) <= (others => '0') ;
	block3x3(2)(2) <= (others => '0') ;
	line_wr <= '0' ;
	k02 <= (others => '0') ;
	k12 <= (others => '0') ;
	pixel_counter <= (others => '0') ;
	pixel_state <= LOAD_VALUES2 ;
elsif clk'event and clk = '1' then
	case pixel_state is
		when LOAD_VALUES1 => -- load value from fifos into buffer
			new_block <= '0' ;
			line_wr <= '0' ;
			pixel_counter <= (pixel_counter + 1) ;
			pixel_state <= LOAD_VALUES2 ;
		when LOAD_VALUES2  =>
			new_block <= '0' ;
			line_wr <= '0' ;
			if nb_line > 0 then
				k12 <= signed('0' & LINE2_OUTPUT) ;
				k02 <= signed('0' & LINE1_OUTPUT) ;
				if hsync = '1' then
					pixel_state <= END_HSYNC ;
				else
					pixel_state <= END_PIXEL ;
				end if ;
			else 
				k12 <= (others => '0') ;
				k02 <= (others => '0') ;
				if hsync = '1' then
						pixel_state <= END_HSYNC ;
				else
					pixel_state <= END_PIXEL ;
				end if ;
			end if;
		when WAIT_PIXEL =>
			new_block <= '0' ;
			line_wr <= '0' ;
			if pixel_clock = '1' and hsync = '0' and vsync = '0' then
				block3x3(0)(2) <= k02 ;
				block3x3(0)(1) <= block3x3(0)(2) ; -- shifting matrix to right
				block3x3(0)(0) <= block3x3(0)(1) ;
				
				block3x3(1)(2) <= k12 ;
				block3x3(1)(1) <= block3x3(1)(2) ;
				block3x3(1)(0) <= block3x3(1)(1) ;
				
				block3x3(2)(2) <= signed('0' & pixel_data_in) ;
				block3x3(2)(1) <= block3x3(2)(2) ;
				block3x3(2)(0) <= block3x3(2)(1) ;
				
				LINE1_input <= std_logic_vector(k12(7 downto 0)) ; -- shifting pixel to upper line fifo
				LINE2_input <= pixel_data_in ; -- shifting pixel to upper line fifo
				line_wr <= '1' ;
				
				new_block <= '1' ;
				pixel_state <= LOAD_VALUES1 ;
			elsif  hsync = '1' then
				pixel_counter <= (others => '0') ;
				pixel_state <= LOAD_VALUES2 ;
			elsif vsync = '1' then
				pixel_counter <= (others => '0') ;
				block3x3(0)(0) <= (others => '0') ;
				block3x3(0)(1) <= (others => '0') ; -- zeroing matrix
				block3x3(0)(2) <= (others => '0') ;
	
				block3x3(1)(0) <= (others => '0') ;
				block3x3(1)(1) <= (others => '0') ;
				block3x3(1)(2) <= (others => '0') ;
	
				block3x3(2)(0) <= (others => '0') ;
				block3x3(2)(1) <= (others => '0') ;
				block3x3(2)(2) <= (others => '0') ;
			end if;
		when END_PIXEL => -- waiting for end of pixel
			new_block <= '0' ;
			line_wr <= '0' ;
			if pixel_clock = '0' then
				pixel_state <= WAIT_PIXEL ;
			elsif  hsync = '1' then
				pixel_state <= LOAD_VALUES2 ;
			end if;
		when END_HSYNC => -- waiting for end of pixel
			new_block <= '0' ;
			line_wr <= '0' ;
			if hsync = '0' then
				pixel_state <= WAIT_PIXEL ;
			end if;
		when others =>
			pixel_state <= WAIT_PIXEL ;
	end case ;
end if;
end process;


process(clk, arazb)
begin
if arazb = '0' then 
	nb_line <= (others => '0') ;
	hsync_state0 <= WAIT_HSYNC ;
elsif clk'event and clk = '1'  then
	case hsync_state0 is
		when WAIT_HSYNC =>
			if hsync = '1' then
				if nb_line < 3 then
					nb_line <= nb_line + 1 ;
				end if;
				hsync_state0 <= END_HSYNC ;
			end if ;
		when END_HSYNC =>
			if vsync = '1' then
				nb_line <= (others => '0') ;
			elsif hsync = '0' then
				hsync_state0 <= WAIT_HSYNC ;
			end if;
		when others =>
			nb_line <= (others => '0') ;
			hsync_state0 <= WAIT_HSYNC ;
	end case ;
end if;
end process;


block_out(0)(2) <= block3x3(0)(2) ;
block_out(1)(2) <= block3x3(1)(2) ;
block_out(2)(2) <= block3x3(2)(2) ;

block_out(0)(1) <= block3x3(0)(1) when pixel_counter > 1 else (others => '0'); -- edges
block_out(1)(1) <= block3x3(1)(1) when pixel_counter > 1 else (others => '0'); -- edges
block_out(2)(1) <= block3x3(2)(1) when pixel_counter > 1 else (others => '0'); -- edges

block_out(0)(0) <= block3x3(0)(0) when pixel_counter > 2 else (others => '0'); -- edges
block_out(1)(0) <= block3x3(1)(0) when pixel_counter > 2 else (others => '0'); -- edges
block_out(2)(0) <= block3x3(2)(0) when pixel_counter > 2 else (others => '0'); -- edges

end Behavioral;

